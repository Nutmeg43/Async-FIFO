package fifo_pkg;
    `include "uvm.sv"
    import uvm_pkg::*;
    `include "fifo_intf.sv"
    `include "fifo_seq.sv"
    `include "fifo_sequence.sv"
    `include "fifo_scoreboard.sv"
    `include "fifo_driver.sv"
    `include "fifo_monitor.sv"
    `include "fifo_agent.sv"
    `include "fifo_env.sv"
    `include "fifo_test.sv"   
endpackage
